module test (input A, output B);
    assign B = A;
endmodule 